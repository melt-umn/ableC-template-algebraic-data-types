grammar edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes;

exports edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:datatype;
exports edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:allocation;