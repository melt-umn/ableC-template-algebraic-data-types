grammar edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:allocation;

exports edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:allocation:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:allocation:concretesyntax;
