grammar edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:datatype;

exports edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:datatype:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:datatype:concretesyntax;
